`timescale 1ns / 1ps

module ALU(
	input clk
);

endmodule
